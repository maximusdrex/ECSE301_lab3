*
* .CONNECT statements
*
.CONNECT GND 0


* ELDO netlist generated with ICnet by 'max' on Mon Mar 21 2022 at 14:05:01

*
* Globals.
*
.global VDD GND

*
* Component pathname : $ADK/parts/inv02
*
.subckt INV02  A Y

        M_I$6 Y A VDD VDD p L=0.6u W=5.4u
        M_I$5 Y A GND GND n L=0.6u W=3u
.ends INV02

*
* Component pathname : $ADK/parts/aoi22
*
.subckt AOI22  B1 A0 A1 B0 Y

        M_I$425 Y B0 N$9 GND n L=0.6u W=3u
        M_I$426 Y B1 N$4 VDD p L=0.6u W=3.9u
        M_I$12 N$8 A1 GND GND n L=0.6u W=3u
        M_I$11 Y A0 N$8 GND n L=0.6u W=3u
        M_I$7 Y B0 N$4 VDD p L=0.6u W=3.9u
        M_I$6 N$4 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$4 A0 VDD VDD p L=0.6u W=3.9u
        M_I$13 N$9 B1 GND GND n L=0.6u W=3u
.ends AOI22

*
* Component pathname : $ADK/parts/xnor2
*
.subckt XNOR2  Y A0 A1

        M_I$218 N$213 A1 GND GND n L=0.6u W=3u
        M_I$217 N$212 A0 N$213 GND n L=0.6u W=3u
        M_I$9 N$212 A1 VDD VDD p L=0.6u W=3.9u
        M_I$8 N$212 A0 VDD VDD p L=0.6u W=3.9u
        M_I$7 N$3 N$212 GND GND n L=0.6u W=3u
        M_I$6 Y A1 N$3 GND n L=0.6u W=3u
        M_I$5 Y A0 N$3 GND n L=0.6u W=3u
        M_I$4 Y A1 N$1 VDD p L=0.6u W=7.8u
        M_I$3 Y N$212 VDD VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends XNOR2

*
* Component pathname : $ADK/parts/mux21_ni
*
.subckt MUX21_NI  S0 A0 A1 Y

        M_I$18 Y N$11 GND GND n L=0.6u W=1.5u
        M_I$17 Y N$11 VDD VDD p L=0.6u W=2.7u
        M_I$16 N$11 S0 N$7 VDD p L=0.6u W=5.4u
        M_I$11 N$3 A1 GND GND n L=0.6u W=3u
        M_I$10 N$11 S0 N$3 GND n L=0.6u W=3u
        M_I$9 N$11 N$4 N$2 VDD p L=0.6u W=5.4u
        M_I$8 N$2 A1 VDD VDD p L=0.6u W=5.4u
        M_I$7 N$1 A0 GND GND n L=0.6u W=3u
        M_I$6 N$11 N$4 N$1 GND n L=0.6u W=3u
        M_I$4 N$7 A0 VDD VDD p L=0.6u W=5.4u
        M_I$3 N$4 S0 GND GND n L=0.6u W=1.5u
        M_I$2 N$4 S0 VDD VDD p L=0.6u W=2.7u
.ends MUX21_NI

*
* Component pathname : $ADK/parts/xor2
*
.subckt XOR2  Y A0 A1

        M_I$421 Y N$4 GND GND n L=0.6u W=1.5u
        M_I$420 Y N$4 VDD VDD p L=0.6u W=2.7u
        M_I$218 N$213 A1 GND GND n L=0.6u W=3u
        M_I$217 N$212 A0 N$213 GND n L=0.6u W=3u
        M_I$9 N$212 A1 VDD VDD p L=0.6u W=3.9u
        M_I$8 N$212 A0 VDD VDD p L=0.6u W=3.9u
        M_I$7 N$3 N$212 GND GND n L=0.6u W=3u
        M_I$6 N$4 A1 N$3 GND n L=0.6u W=3u
        M_I$5 N$4 A0 N$3 GND n L=0.6u W=3u
        M_I$4 N$4 A1 N$1 VDD p L=0.6u W=7.8u
        M_I$3 N$4 N$212 VDD VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends XOR2

*
* Component pathname : /home/max/301/ECSE301_lab3/AddSub_S/AddSub
*
.subckt ADDSUB  MULT[0] MULT[1] MULT[2] MULT[3] A_IN[0] A_IN[1] A_IN[2]
+ A_IN[3] A_OUT[0] A_OUT[1] A_OUT[2] A_OUT[3] CLOCK CONTROL

        X_IX213 NX10 NX212 INV02
        X_IX211 NX12 NX212 A_IN[1] NX32 NX210 AOI22
        X_IX43 NX42 MULT[3] CONTROL XNOR2
        X_IX45 NX44 A_IN[3] NX42 XNOR2
        X_IX47 A_OUT[3] NX219 NX44 XNOR2
        X_IX1 NX0 MULT[2] CONTROL XNOR2
        X_IX3 NX2 A_IN[2] NX0 XNOR2
        X_IX49 A_OUT[2] NX210 NX2 XNOR2
        X_IX11 NX10 MULT[1] CONTROL XNOR2
        X_IX13 NX12 A_IN[1] NX10 XNOR2
        X_IX220 NX2 NX0 NX210 NX219 MUX21_NI
        X_IX33 MULT[0] CONTROL A_IN[0] NX32 MUX21_NI
        X_IX51 A_OUT[1] NX32 NX12 XOR2
        X_IX53 A_OUT[0] A_IN[0] MULT[0] XOR2
.ends ADDSUB

*
* Component pathname : $ADK/parts/nand02_2x
*
.subckt NAND02_2X  Y A0 A1

        M_I$9 Y A1 VDD VDD p L=0.6u W=6u
        M_I$8 Y A0 VDD VDD p L=0.6u W=6u
        M_I$3 Y A0 N$5 GND n L=0.6u W=6u
        M_I$2 N$5 A1 GND GND n L=0.6u W=6u
.ends NAND02_2X

*
* Component pathname : $ADK/parts/nor02_2x
*
.subckt NOR02_2X  A0 A1 Y

        M_I$5 Y A0 GND GND n L=0.6u W=3u
        M_I$4 Y A1 GND GND n L=0.6u W=3u
        M_I$3 Y A1 N$1 VDD p L=0.6u W=7.8u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends NOR02_2X

*
* Component pathname : $ADK/parts/ao22
*
.subckt AO22  A1 A0 B0 Y B1

        M_I$16 Y N$215 VDD VDD p L=0.6u W=2.7u
        M_I$18 Y N$215 GND GND n L=0.6u W=1.5u
        M_I$14 N$215 B0 N$2 GND n L=0.6u W=3u
        M_I$13 N$215 B1 N$6 VDD p L=0.6u W=3.9u
        M_I$12 N$1 A1 GND GND n L=0.6u W=3u
        M_I$11 N$215 A0 N$1 GND n L=0.6u W=3u
        M_I$7 N$215 B0 N$6 VDD p L=0.6u W=3.9u
        M_I$6 N$6 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$6 A0 VDD VDD p L=0.6u W=3.9u
        M_I$4 N$2 B1 GND GND n L=0.6u W=3u
.ends AO22

*
* Component pathname : $ADK/parts/ao32
*
.subckt AO32  Y A0 A1 A2 B0 B1

        M_I$222 Y N$214 GND GND n L=0.6u W=1.5u
        M_I$221 Y N$214 VDD VDD p L=0.6u W=2.7u
        M_I$12 N$6 B1 GND GND n L=0.6u W=3u
        M_I$11 N$214 B0 N$6 GND n L=0.6u W=3u
        M_I$10 N$5 A2 GND GND n L=0.6u W=4.5u
        M_I$9 N$4 A1 N$5 GND n L=0.6u W=4.5u
        M_I$8 N$214 A0 N$4 GND n L=0.6u W=4.5u
        M_I$6 N$214 B0 N$11 VDD p L=0.6u W=3.9u
        M_I$5 N$214 B1 N$11 VDD p L=0.6u W=3.9u
        M_I$4 N$11 A0 VDD VDD p L=0.6u W=3.9u
        M_I$3 N$11 A1 VDD VDD p L=0.6u W=3.9u
        M_I$2 N$11 A2 VDD VDD p L=0.6u W=3.9u
.ends AO32

*
* Component pathname : $ADK/parts/dff
*
.subckt DFF  QB Q CLK D

        M_I$441 N$847 BCLK- N$851 GND n L=0.6u W=4.5u
        M_I$440 N$849 N$847 VDD VDD p L=0.6u W=1.5u
        M_I$439 N$847 BCLK- N$848 VDD p L=0.6u W=1.5u
        M_I$438 N$848 N$849 VDD VDD p L=0.6u W=1.5u
        M_I$437 N$847 BCLK N$845 VDD p L=0.6u W=8.1u
        M_I$436 N$845 D VDD VDD p L=0.6u W=8.1u
        M_I$452 BCLK BCLK- GND GND n L=0.6u W=3u
        M_I$673 Q QB GND GND n L=0.6u W=3u
        M_I$672 Q QB VDD VDD p L=0.6u W=5.4u
        M_I$669 QB N$1074 GND GND n L=0.6u W=3u
        M_I$675 QB N$1074 VDD VDD p L=0.6u W=5.4u
        M_I$668 N$1071 N$1074 GND GND n L=0.6u W=1.5u
        M_I$667 N$1073 N$1071 GND GND n L=0.6u W=1.5u
        M_I$666 N$1074 BCLK- N$1073 GND n L=0.6u W=1.5u
        M_I$665 N$1072 N$847 GND GND n L=0.6u W=4.5u
        M_I$664 N$1074 BCLK N$1072 GND n L=0.6u W=4.5u
        M_I$663 N$1071 N$1074 VDD VDD p L=0.6u W=1.5u
        M_I$662 N$1074 BCLK N$1070 VDD p L=0.6u W=1.5u
        M_I$661 N$1070 N$1071 VDD VDD p L=0.6u W=1.5u
        M_I$660 N$1074 BCLK- N$1069 VDD p L=0.6u W=8.1u
        M_I$659 N$1069 N$847 VDD VDD p L=0.6u W=8.1u
        M_I$449 BCLK- CLK GND GND n L=0.6u W=3u
        M_I$448 BCLK- CLK VDD VDD p L=0.6u W=5.4u
        M_I$453 BCLK BCLK- VDD VDD p L=0.6u W=5.4u
        M_I$445 N$849 N$847 GND GND n L=0.6u W=1.5u
        M_I$444 N$852 N$849 GND GND n L=0.6u W=1.5u
        M_I$443 N$847 BCLK N$852 GND n L=0.6u W=1.5u
        M_I$442 N$851 D GND GND n L=0.6u W=4.5u
.ends DFF

*
* Component pathname : /home/max/301/ECSE301_lab3/Qreg_S/Qreg
*
.subckt QREG  LOAD[0] LOAD[1] LOAD[2] LOAD[3] CONTROL[0] CONTROL[1] Q_OUT[0]
+ Q_OUT[1] Q_OUT[2] Q_OUT[3] Q_OUT[4] A_IN CLOCK

        X_IX209 NX4 NX208 INV02
        X_IX207 CONTROL[0] NX206 INV02
        X_IX201 CLOCK NOT_CLOCK INV02
        X_IX5 NX4 CONTROL[1] CONTROL[0] NAND02_2X
        X_IX11 CONTROL[0] CONTROL[1] NX10 NOR02_2X
        X_IX23 CONTROL[1] A_IN LOAD[3] NX22 NX10 AO22
        X_IX35 Q_OUT[4] CONTROL[1] LOAD[2] NX34 NX10 AO22
        X_IX45 Q_OUT[3] CONTROL[1] LOAD[1] NX44 NX10 AO22
        X_IX55 Q_OUT[2] CONTROL[1] LOAD[0] NX54 NX10 AO22
        X_IX135 NX4 Q_OUT[4] NX22 NX134 MUX21_NI
        X_IX145 NX4 Q_OUT[3] NX34 NX144 MUX21_NI
        X_IX155 NX4 Q_OUT[2] NX44 NX154 MUX21_NI
        X_IX165 NX4 Q_OUT[1] NX54 NX164 MUX21_NI
        X_IX175 NX174 CONTROL[1] Q_OUT[1] NX206 Q_OUT[0] NX208 AO32
        X_REG_Q_OUT_4 N$DUMMY_ESC1[4] Q_OUT[4] NOT_CLOCK NX134 DFF
        X_REG_Q_OUT_3 N$DUMMY_ESC1[3] Q_OUT[3] NOT_CLOCK NX144 DFF
        X_REG_Q_OUT_2 N$DUMMY_ESC1[2] Q_OUT[2] NOT_CLOCK NX154 DFF
        X_REG_Q_OUT_1 N$DUMMY_ESC1[1] Q_OUT[1] NOT_CLOCK NX164 DFF
        X_REG_Q_OUT_0 N$DUMMY_ESC1[0] Q_OUT[0] NOT_CLOCK NX174 DFF
.ends QREG

*
* Component pathname : $ADK/parts/nor03
*
.subckt NOR03  A2 A0 A1 Y

        M_I$213 Y A0 GND GND n L=0.6u W=1.8u
        M_I$211 Y A2 N$211 VDD p L=0.6u W=8.1u
        M_I$5 Y A1 GND GND n L=0.6u W=1.8u
        M_I$4 Y A2 GND GND n L=0.6u W=1.8u
        M_I$3 N$211 A1 N$1 VDD p L=0.6u W=8.1u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=8.1u
.ends NOR03

*
* Component pathname : $ADK/parts/ao21
*
.subckt AO21  A1 A0 B0 Y

        M_I$14 Y N$3 VDD VDD p L=0.6u W=2.7u
        M_I$13 Y N$3 GND GND n L=0.6u W=1.5u
        M_I$12 N$2 A1 GND GND n L=0.6u W=3u
        M_I$11 N$3 A0 N$2 GND n L=0.6u W=3u
        M_I$7 N$3 B0 N$1 VDD p L=0.6u W=3.9u
        M_I$6 N$1 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$1 A0 VDD VDD p L=0.6u W=3.9u
        M_I$4 N$3 B0 GND GND n L=0.6u W=1.5u
.ends AO21

*
* Component pathname : /home/max/301/ECSE301_lab3/Areg_S/Areg
*
.subckt AREG  ADDER[0] ADDER[1] ADDER[2] ADDER[3] CONTROL[0] CONTROL[1]
+ A_OUT[0] A_OUT[1] A_OUT[2] A_OUT[3] CLOCK

        X_IX5 NX4 CONTROL[1] CONTROL[0] NAND02_2X
        X_IX11 CONTROL[0] CONTROL[1] NX10 NOR02_2X
        X_IX164 ADDER[3] NX163 INV02
        X_IX110 CONTROL[1] NX163 CONTROL[0] NX109 NOR03
        X_IX112 CONTROL[1] A_OUT[3] NX109 NX111 AO21
        X_IX33 A_OUT[3] CONTROL[1] ADDER[2] NX32 NX10 AO22
        X_IX43 A_OUT[2] CONTROL[1] ADDER[1] NX42 NX10 AO22
        X_IX53 A_OUT[1] CONTROL[1] ADDER[0] NX52 NX10 AO22
        X_IX122 NX4 A_OUT[2] NX32 NX121 MUX21_NI
        X_IX132 NX4 A_OUT[1] NX42 NX131 MUX21_NI
        X_IX142 NX4 A_OUT[0] NX52 NX141 MUX21_NI
        X_REG_A_OUT_3 N$DUMMY_ESC1[3] A_OUT[3] CLOCK NX111 DFF
        X_REG_A_OUT_2 N$DUMMY_ESC1[2] A_OUT[2] CLOCK NX121 DFF
        X_REG_A_OUT_1 N$DUMMY_ESC1[1] A_OUT[1] CLOCK NX131 DFF
        X_REG_A_OUT_0 N$DUMMY_ESC1[0] A_OUT[0] CLOCK NX141 DFF
.ends AREG

*
* Component pathname : /home/max/301/ECSE301_lab3/Mreg_S/Mreg
*
.subckt MREG  LOAD[0] LOAD[1] LOAD[2] LOAD[3] M_OUT[0] M_OUT[1] M_OUT[2]
+ M_OUT[3] CLOCK CONTROL

        X_IX152 CONTROL M_OUT[3] LOAD[3] NX151 MUX21_NI
        X_IX142 CONTROL M_OUT[2] LOAD[2] NX141 MUX21_NI
        X_IX132 CONTROL M_OUT[1] LOAD[1] NX131 MUX21_NI
        X_IX122 CONTROL M_OUT[0] LOAD[0] NX121 MUX21_NI
        X_REG_M_OUT_3 N$DUMMY_ESC1[3] M_OUT[3] CLOCK NX151 DFF
        X_REG_M_OUT_2 N$DUMMY_ESC1[2] M_OUT[2] CLOCK NX141 DFF
        X_REG_M_OUT_1 N$DUMMY_ESC1[1] M_OUT[1] CLOCK NX131 DFF
        X_REG_M_OUT_0 N$DUMMY_ESC1[0] M_OUT[0] CLOCK NX121 DFF
.ends MREG

*
* Component pathname : $ADK/parts/nor02ii
*
.subckt NOR02II  A0 A1 Y

        MP1 N$208 A1 VDD VDD p L=0.6u W=2.7u
        MN1 N$208 A1 GND GND n L=0.6u W=1.5u
        MN4 Y A0 GND GND n L=0.6u W=1.5u
        MN2 Y N$208 GND GND n L=0.6u W=1.5u
        MP4 Y N$208 N$4 VDD p L=0.6u W=3.9u
        MP2 N$4 A0 VDD VDD p L=0.6u W=3.9u
.ends NOR02II

*
* Component pathname : $ADK/parts/latch
*
.subckt LATCH  Q CLK D

        M_I$222 Q N$17 GND GND n L=0.6u W=1.5u
        M_I$221 Q N$17 VDD VDD p L=0.6u W=2.7u
        M_I$15 N$10 CLK GND GND n L=0.6u W=1.5u
        M_I$13 N$222 N$17 GND GND n L=0.6u W=1.5u
        M_I$12 N$15 N$222 GND GND n L=0.6u W=1.5u
        M_I$11 N$17 N$10 N$15 GND n L=0.6u W=1.5u
        M_I$10 N$13 D GND GND n L=0.6u W=4.5u
        M_I$9 N$17 CLK N$13 GND n L=0.6u W=4.5u
        M_I$6 N$17 CLK N$15 VDD p L=0.6u W=1.5u
        M_I$7 N$222 N$17 VDD VDD p L=0.6u W=2.7u
        M_I$5 N$15 N$222 VDD VDD p L=0.6u W=1.5u
        M_I$4 N$17 N$10 N$11 VDD p L=0.6u W=8.1u
        M_I$3 N$11 D VDD VDD p L=0.6u W=8.1u
        M_I$2 N$10 CLK VDD VDD p L=0.6u W=2.7u
.ends LATCH

*
* Component pathname : $ADK/parts/and02
*
.subckt AND02  Y A0 A1

        M_I$674 Y N$5 VDD VDD p L=0.6u W=2.7u
        M_I$675 Y N$5 GND GND n L=0.6u W=1.5u
        M_I$472 N$5 A1 VDD VDD p L=0.6u W=3.6u
        M_I$471 N$5 A0 VDD VDD p L=0.6u W=3.6u
        M_I$4 N$5 A0 N$7 GND n L=0.6u W=3u
        M_I$5 N$7 A1 GND GND n L=0.6u W=3u
.ends AND02

*
* Component pathname : $ADK/parts/oai21
*
.subckt OAI21  A0 A1 B0 Y

        M_I$5 N$7 B0 GND GND n L=0.6u W=3u
        M_I$4 Y A1 N$7 GND n L=0.6u W=3u
        M_I$3 Y A0 N$7 GND n L=0.6u W=3u
        M_I$12 Y B0 VDD VDD p L=0.6u W=3.6u
        M_I$2 Y A1 N$9 VDD p L=0.6u W=7.2u
        M_I$1 N$9 A0 VDD VDD p L=0.6u W=7.2u
.ends OAI21

*
* Component pathname : $ADK/parts/inv01
*
.subckt INV01  A Y

        M_I$411 Y A VDD VDD p L=0.6u W=2.7u
        M_I$412 Y A GND GND n L=0.6u W=1.5u
.ends INV01

*
* Component pathname : $ADK/parts/latchr
*
.subckt LATCHR  QB R CLK D

        M_I$1954 N$3723 R GND GND n L=0.6u W=3u
        M_I$1953 N$3723 R N$3722 VDD p L=0.6u W=3.6u
        M_I$1244 N$3516 N$3723 VDD VDD p L=0.6u W=1.5u
        M_I$1245 N$3108 N$3723 GND GND n L=0.6u W=1.5u
        M_I$1749 N$3723 N$3929 GND GND n L=0.6u W=3u
        M_I$1240 N$3929 CLK N$3516 VDD p L=0.6u W=1.5u
        M_I$15 N$3100 CLK GND GND n L=0.6u W=1.5u
        M_I$1242 N$3722 N$3929 VDD VDD p L=0.6u W=3.6u
        M_I$1036 QB N$3723 GND GND n L=0.6u W=1.5u
        M_I$10 N$13 D GND GND n L=0.6u W=4.5u
        M_I$9 N$3929 CLK N$13 GND n L=0.6u W=4.5u
        M_I$1035 QB N$3723 VDD VDD p L=0.6u W=2.7u
        M_I$1447 N$3929 N$3100 N$3108 GND n L=0.6u W=1.5u
        M_I$4 N$3929 N$3100 N$11 VDD p L=0.6u W=8.1u
        M_I$3 N$11 D VDD VDD p L=0.6u W=8.1u
        M_I$2 N$3100 CLK VDD VDD p L=0.6u W=2.7u
.ends LATCHR

*
* Component pathname : $ADK/parts/or03
*
.subckt OR03  A2 A0 A1 Y

        M_I$416 Y N$214 GND GND n L=0.6u W=1.5u
        M_I$415 Y N$214 VDD VDD p L=0.6u W=2.7u
        M_I$213 N$214 A0 GND GND n L=0.6u W=1.8u
        M_I$211 N$214 A2 N$211 VDD p L=0.6u W=8.1u
        M_I$5 N$214 A1 GND GND n L=0.6u W=1.8u
        M_I$4 N$214 A2 GND GND n L=0.6u W=1.8u
        M_I$3 N$211 A1 N$1 VDD p L=0.6u W=8.1u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=8.1u
.ends OR03

*
* Component pathname : $ADK/parts/buf08
*
.subckt BUF08  A Y

        M_I$1023 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$1022 Y N$411 GND GND n L=0.6u W=3u
        M_I$1021 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$1020 Y N$411 GND GND n L=0.6u W=3u
        M_I$817 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$818 Y N$411 GND GND n L=0.6u W=3u
        M_I$614 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$615 Y N$411 GND GND n L=0.6u W=3u
        M_I$411 N$411 A VDD VDD p L=0.6u W=5.4u
        M_I$412 N$411 A GND GND n L=0.6u W=3u
.ends BUF08

*
* Component pathname : $ADK/parts/buf02
*
.subckt BUF02  A Y

        M_I$614 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$615 Y N$411 GND GND n L=0.6u W=3u
        M_I$411 N$411 A VDD VDD p L=0.6u W=2.7u
        M_I$412 N$411 A GND GND n L=0.6u W=1.5u
.ends BUF02

*
* Component pathname : $ADK/parts/inv08
*
.subckt INV08  A Y

        M_I$618 Y A GND GND n L=0.6u W=3u
        M_I$617 Y A VDD VDD p L=0.6u W=5.4u
        M_I$616 Y A GND GND n L=0.6u W=3u
        M_I$619 Y A VDD VDD p L=0.6u W=5.4u
        M_I$412 Y A VDD VDD p L=0.6u W=5.4u
        M_I$413 Y A GND GND n L=0.6u W=3u
        M_I$6 Y A VDD VDD p L=0.6u W=5.4u
        M_I$5 Y A GND GND n L=0.6u W=3u
.ends INV08

*
* Component pathname : $ADK/parts/nor03_2x
*
.subckt NOR03_2X  A1 A0 A2 Y

        M_I$12 Y A0 GND GND n L=0.6u W=3.3u
        M_I$10 Y A2 N$3 VDD p L=0.6u W=12u
        M_I$5 Y A1 GND GND n L=0.6u W=3.3u
        M_I$4 Y A2 GND GND n L=0.6u W=3.3u
        M_I$3 N$3 A1 N$1 VDD p L=0.6u W=12u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=12u
.ends NOR03_2X

*
* Component pathname : $ADK/parts/nor04
*
.subckt NOR04  A3 A2 A0 A1 Y

        M_I$415 Y A3 GND GND n L=0.6u W=3u
        M_I$416 Y A3 N$418 VDD p L=0.6u W=10.8u
        M_I$213 Y A0 GND GND n L=0.6u W=3u
        M_I$211 N$418 A2 N$211 VDD p L=0.6u W=10.8u
        M_I$5 Y A1 GND GND n L=0.6u W=3u
        M_I$4 Y A2 GND GND n L=0.6u W=3u
        M_I$3 N$211 A1 N$1 VDD p L=0.6u W=10.8u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=10.8u
.ends NOR04

*
* Component pathname : $ADK/parts/or02
*
.subckt OR02  A0 A1 Y

        M_I$212 Y N$5 GND GND n L=0.6u W=1.5u
        M_I$211 Y N$5 VDD VDD p L=0.6u W=2.7u
        M_I$5 N$5 A0 GND GND n L=0.6u W=1.5u
        M_I$4 N$5 A1 GND GND n L=0.6u W=1.5u
        M_I$3 N$5 A1 N$1 VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=3.9u
.ends OR02

*
* Component pathname : /home/max/301/ECSE301_lab3/Control_S/ControlLogic
*
.subckt CONTROLLOGIC  Q_IN[0] Q_IN[1] Q_SIG[0] Q_SIG[1] A_SIG[0] A_SIG[1]
+ ADDER_SIG M_SIG DONE_SIG START CLOCK

        X_IX593 PRES_STATE_0 PRES_STATE_4 PRES_STATE_5 NX592 NOR03
        X_IX5 NX587 NX569 Q_IN[1] NX4 NOR03
        X_IX191 Q_IN[0] NX569 NX630 NX190 NOR03
        X_IX91 NX574 NX622 NX90 NOR02II
        X_IX610 COUNT_1 NX622 NX609 NOR02II
        X_IX141 START NEXT_STATE_5 NX140 NOR02II
        X_IX47 START NEXT_STATE_1 NX46 NOR02II
        X_IX73 START NEXT_STATE_3 NX72 NOR02II
        X_IX179 START NEXT_STATE_0 NX178 NOR02II
        X_IX201 START NEXT_STATE_2 NX200 NOR02II
        X_REG_PRES_STATE_3 NX574 PRES_STATE_3 CLOCK NX72 DFF
        X_REG_PRES_STATE_4 NOT_PRES_STATE_4 PRES_STATE_4 CLOCK NX158 DFF
        X_REG_PRES_STATE_5 NX598 PRES_STATE_5 CLOCK NX140 DFF
        X_REG_PRES_STATE_1 N$DUMMY_ESC1[1] PRES_STATE_1 CLOCK NX46 DFF
        X_REG_PRES_STATE_0 NX569 PRES_STATE_0 CLOCK NX178 DFF
        X_REG_PRES_STATE_2 N$DUMMY_ESC1[0] PRES_STATE_2 CLOCK NX200 DFF
        X_LAT_Q_SIG_1 Q_SIG[1] NX648 NOT_PRES_STATE_4 LATCH
        X_LAT_Q_SIG_0 Q_SIG[0] NX648 NX10 LATCH
        X_LAT_A_SIG_1 A_SIG[1] NX648 NX24 LATCH
        X_LAT_A_SIG_0 A_SIG[0] NX648 NX28 LATCH
        X_LAT_DONE_SIG DONE_SIG NX648 PRES_STATE_5 LATCH
        X_LAT_M_SIG M_SIG NX648 PRES_STATE_4 LATCH
        X_LAT_COUNT_1 COUNT_1 NX14 NX80 LATCH
        X_LAT_COUNT_2 COUNT_2 NX14 NX108 LATCH
        X_LAT_NEXT_STATE_5 NEXT_STATE_5 NX646 NX130 LATCH
        X_LAT_NEXT_STATE_4 NEXT_STATE_4 NX646 NX150 LATCH
        X_LAT_NEXT_STATE_1 NEXT_STATE_1 NX646 NX4 LATCH
        X_LAT_NEXT_STATE_3 NEXT_STATE_3 NX646 NX62 LATCH
        X_LAT_NEXT_STATE_0 NEXT_STATE_0 NX646 NX168 LATCH
        X_LAT_NEXT_STATE_2 NEXT_STATE_2 NX646 NX190 LATCH
        X_LAT_ADDER_SIG ADDER_SIG NX646 PRES_STATE_2 LATCH
        X_IX81 NX80 PRES_STATE_3 NX556 AND02
        X_IX626 PRES_STATE_4 PRES_STATE_3 CLOCK NX625 OAI21
        X_IX109 NX574 NX607 NOT_PRES_STATE_4 NX108 OAI21
        X_IX11 PRES_STATE_4 PRES_STATE_3 NX10 NOR02_2X
        X_IX151 START NX598 NX150 NOR02_2X
        X_LAT_COUNT_0__U2 NX5 COUNT_0 INV01
        X_LAT_COUNT_0__U1 NX5 GND NX14 NX650 LATCHR
        X_IX629 COUNT_1 COUNT_2 NX622 NX656 OR03
        X_IX649 NX90 NX650 BUF08
        X_IX660 NX609 NX661 BUF02
        X_LAT_COUNT_0__U3 NX5 NX622 BUF02
        X_IX647 NX36 NX648 BUF02
        X_IX645 NX36 NX646 BUF02
        X_IX15 NX625 NX14 INV08
        X_IX25 PRES_STATE_4 PRES_STATE_1 PRES_STATE_2 NX24 NOR03_2X
        X_IX127 COUNT_1 NX622 NX574 COUNT_2 NX126 NOR04
        X_IX37 NX36 NX590 NX625 NAND02_2X
        X_IX29 NX592 NX28 INV02
        X_IX631 Q_IN[1] NX630 INV02
        X_IX617 CLOCK NX616 INV02
        X_IX588 Q_IN[0] NX587 INV02
        X_IX608 NX607 COUNT_2 NX661 XNOR2
        X_IX582 NX581 Q_IN[1] Q_IN[0] XNOR2
        X_IX169 NX656 PRES_STATE_3 PRES_STATE_4 NX168 AO21
        X_IX105 COUNT_0 COUNT_1 NX661 NX556 AO21
        X_IX131 PRES_STATE_5 START NX126 NX130 AO21
        X_IX591 NX24 NX592 NX616 NX590 AO21
        X_IX61 NX581 PRES_STATE_0 PRES_STATE_1 NX60 AO21
        X_IX159 NEXT_STATE_4 START NX158 OR02
        X_IX63 NX60 PRES_STATE_2 NX62 OR02
.ends CONTROLLOGIC

*
* MAIN CELL: Component pathname : /home/max/301/ECSE301_lab3/TopModel
*
        X_ADDSUB1 MULT[0] MULT[1] MULT[2] MULT[3] OUT[4] OUT[5] OUT[6] OUT[7]
+ ADDER[0] ADDER[1] ADDER[2] ADDER[3] CLK N$31 ADDSUB
        X_QREG1 Q_IN[0] Q_IN[1] Q_IN[2] Q_IN[3] Q_SIG[0] Q_SIG[1] Q_OUT[0]
+ OUT[0] OUT[1] OUT[2] OUT[3] OUT[4] CLK QREG
        X_AREG1 ADDER[0] ADDER[1] ADDER[2] ADDER[3] A_SIG[0] A_SIG[1] OUT[4]
+ OUT[5] OUT[6] OUT[7] CLK AREG
        X_MREG1 M_IN[0] M_IN[1] M_IN[2] M_IN[3] MULT[0] MULT[1] MULT[2]
+ MULT[3] CLK N$33 MREG
        X_CONTROLLOGIC1 Q_OUT[0] OUT[0] Q_SIG[0] Q_SIG[1] A_SIG[0] A_SIG[1]
+ N$31 N$33 DONE START CLK CONTROLLOGIC
*
.end
