*
* .CONNECT statements
*
.CONNECT GND 0


* ELDO netlist generated with ICnet by 'max' on Thu Mar  3 2022 at 13:35:32

*
* Globals.
*
.global VDD GND

*
* Component pathname : $ADK/parts/inv02
*
.subckt INV02  A Y

        M_I$6 Y A VDD VDD p L=0.6u W=5.4u
        M_I$5 Y A GND GND n L=0.6u W=3u
.ends INV02

*
* Component pathname : $ADK/parts/aoi22
*
.subckt AOI22  B1 A0 A1 B0 Y

        M_I$425 Y B0 N$9 GND n L=0.6u W=3u
        M_I$426 Y B1 N$4 VDD p L=0.6u W=3.9u
        M_I$12 N$8 A1 GND GND n L=0.6u W=3u
        M_I$11 Y A0 N$8 GND n L=0.6u W=3u
        M_I$7 Y B0 N$4 VDD p L=0.6u W=3.9u
        M_I$6 N$4 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$4 A0 VDD VDD p L=0.6u W=3.9u
        M_I$13 N$9 B1 GND GND n L=0.6u W=3u
.ends AOI22

*
* Component pathname : $ADK/parts/xnor2
*
.subckt XNOR2  Y A0 A1

        M_I$218 N$213 A1 GND GND n L=0.6u W=3u
        M_I$217 N$212 A0 N$213 GND n L=0.6u W=3u
        M_I$9 N$212 A1 VDD VDD p L=0.6u W=3.9u
        M_I$8 N$212 A0 VDD VDD p L=0.6u W=3.9u
        M_I$7 N$3 N$212 GND GND n L=0.6u W=3u
        M_I$6 Y A1 N$3 GND n L=0.6u W=3u
        M_I$5 Y A0 N$3 GND n L=0.6u W=3u
        M_I$4 Y A1 N$1 VDD p L=0.6u W=7.8u
        M_I$3 Y N$212 VDD VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends XNOR2

*
* Component pathname : $ADK/parts/mux21_ni
*
.subckt MUX21_NI  S0 A0 A1 Y

        M_I$18 Y N$11 GND GND n L=0.6u W=1.5u
        M_I$17 Y N$11 VDD VDD p L=0.6u W=2.7u
        M_I$16 N$11 S0 N$7 VDD p L=0.6u W=5.4u
        M_I$11 N$3 A1 GND GND n L=0.6u W=3u
        M_I$10 N$11 S0 N$3 GND n L=0.6u W=3u
        M_I$9 N$11 N$4 N$2 VDD p L=0.6u W=5.4u
        M_I$8 N$2 A1 VDD VDD p L=0.6u W=5.4u
        M_I$7 N$1 A0 GND GND n L=0.6u W=3u
        M_I$6 N$11 N$4 N$1 GND n L=0.6u W=3u
        M_I$4 N$7 A0 VDD VDD p L=0.6u W=5.4u
        M_I$3 N$4 S0 GND GND n L=0.6u W=1.5u
        M_I$2 N$4 S0 VDD VDD p L=0.6u W=2.7u
.ends MUX21_NI

*
* Component pathname : $ADK/parts/xor2
*
.subckt XOR2  Y A0 A1

        M_I$421 Y N$4 GND GND n L=0.6u W=1.5u
        M_I$420 Y N$4 VDD VDD p L=0.6u W=2.7u
        M_I$218 N$213 A1 GND GND n L=0.6u W=3u
        M_I$217 N$212 A0 N$213 GND n L=0.6u W=3u
        M_I$9 N$212 A1 VDD VDD p L=0.6u W=3.9u
        M_I$8 N$212 A0 VDD VDD p L=0.6u W=3.9u
        M_I$7 N$3 N$212 GND GND n L=0.6u W=3u
        M_I$6 N$4 A1 N$3 GND n L=0.6u W=3u
        M_I$5 N$4 A0 N$3 GND n L=0.6u W=3u
        M_I$4 N$4 A1 N$1 VDD p L=0.6u W=7.8u
        M_I$3 N$4 N$212 VDD VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends XOR2

*
* Component pathname : /home/max/EECS301/lab3/AddSub_S/AddSub
*
.subckt ADDSUB  MULT[0] MULT[1] MULT[2] MULT[3] A_IN[0] A_IN[1] A_IN[2]
+ A_IN[3] A_OUT[0] A_OUT[1] A_OUT[2] A_OUT[3] CLOCK CONTROL

        X_IX213 NX10 NX212 INV02
        X_IX211 NX12 NX212 A_IN[1] NX32 NX210 AOI22
        X_IX43 NX42 MULT[3] CONTROL XNOR2
        X_IX45 NX44 A_IN[3] NX42 XNOR2
        X_IX47 A_OUT[3] NX219 NX44 XNOR2
        X_IX1 NX0 MULT[2] CONTROL XNOR2
        X_IX3 NX2 A_IN[2] NX0 XNOR2
        X_IX49 A_OUT[2] NX210 NX2 XNOR2
        X_IX11 NX10 MULT[1] CONTROL XNOR2
        X_IX13 NX12 A_IN[1] NX10 XNOR2
        X_IX220 NX2 NX0 NX210 NX219 MUX21_NI
        X_IX33 MULT[0] CONTROL A_IN[0] NX32 MUX21_NI
        X_IX51 A_OUT[1] NX32 NX12 XOR2
        X_IX53 A_OUT[0] A_IN[0] MULT[0] XOR2
.ends ADDSUB

*
* Component pathname : $ADK/parts/dff
*
.subckt DFF  QB Q CLK D

        M_I$441 N$847 BCLK- N$851 GND n L=0.6u W=4.5u
        M_I$440 N$849 N$847 VDD VDD p L=0.6u W=1.5u
        M_I$439 N$847 BCLK- N$848 VDD p L=0.6u W=1.5u
        M_I$438 N$848 N$849 VDD VDD p L=0.6u W=1.5u
        M_I$437 N$847 BCLK N$845 VDD p L=0.6u W=8.1u
        M_I$436 N$845 D VDD VDD p L=0.6u W=8.1u
        M_I$452 BCLK BCLK- GND GND n L=0.6u W=3u
        M_I$673 Q QB GND GND n L=0.6u W=3u
        M_I$672 Q QB VDD VDD p L=0.6u W=5.4u
        M_I$669 QB N$1074 GND GND n L=0.6u W=3u
        M_I$675 QB N$1074 VDD VDD p L=0.6u W=5.4u
        M_I$668 N$1071 N$1074 GND GND n L=0.6u W=1.5u
        M_I$667 N$1073 N$1071 GND GND n L=0.6u W=1.5u
        M_I$666 N$1074 BCLK- N$1073 GND n L=0.6u W=1.5u
        M_I$665 N$1072 N$847 GND GND n L=0.6u W=4.5u
        M_I$664 N$1074 BCLK N$1072 GND n L=0.6u W=4.5u
        M_I$663 N$1071 N$1074 VDD VDD p L=0.6u W=1.5u
        M_I$662 N$1074 BCLK N$1070 VDD p L=0.6u W=1.5u
        M_I$661 N$1070 N$1071 VDD VDD p L=0.6u W=1.5u
        M_I$660 N$1074 BCLK- N$1069 VDD p L=0.6u W=8.1u
        M_I$659 N$1069 N$847 VDD VDD p L=0.6u W=8.1u
        M_I$449 BCLK- CLK GND GND n L=0.6u W=3u
        M_I$448 BCLK- CLK VDD VDD p L=0.6u W=5.4u
        M_I$453 BCLK BCLK- VDD VDD p L=0.6u W=5.4u
        M_I$445 N$849 N$847 GND GND n L=0.6u W=1.5u
        M_I$444 N$852 N$849 GND GND n L=0.6u W=1.5u
        M_I$443 N$847 BCLK N$852 GND n L=0.6u W=1.5u
        M_I$442 N$851 D GND GND n L=0.6u W=4.5u
.ends DFF

*
* Component pathname : /home/max/EECS301/lab3/Mreg_S/Mreg
*
.subckt MREG  LOAD[0] LOAD[1] LOAD[2] LOAD[3] M_OUT[0] M_OUT[1] M_OUT[2]
+ M_OUT[3] CLOCK CONTROL

        X_IX175 CLOCK NOT_CLOCK INV02
        X_IX162 CONTROL M_3 LOAD[3] NX161 MUX21_NI
        X_IX152 CONTROL M_2 LOAD[2] NX151 MUX21_NI
        X_IX142 CONTROL M_1 LOAD[1] NX141 MUX21_NI
        X_IX132 CONTROL M_0 LOAD[0] NX131 MUX21_NI
        X_REG_M_3 N$DUMMY_ESC1[7] M_3 NOT_CLOCK NX161 DFF
        X_REG_MO_3 N$DUMMY_ESC1[6] M_OUT[3] CLOCK M_3 DFF
        X_REG_M_2 N$DUMMY_ESC1[5] M_2 NOT_CLOCK NX151 DFF
        X_REG_MO_2 N$DUMMY_ESC1[4] M_OUT[2] CLOCK M_2 DFF
        X_REG_M_1 N$DUMMY_ESC1[3] M_1 NOT_CLOCK NX141 DFF
        X_REG_MO_1 N$DUMMY_ESC1[2] M_OUT[1] CLOCK M_1 DFF
        X_REG_M_0 N$DUMMY_ESC1[1] M_0 NOT_CLOCK NX131 DFF
        X_REG_MO_0 N$DUMMY_ESC1[0] M_OUT[0] CLOCK M_0 DFF
.ends MREG

*
* Component pathname : $ADK/parts/nand02_2x
*
.subckt NAND02_2X  Y A0 A1

        M_I$9 Y A1 VDD VDD p L=0.6u W=6u
        M_I$8 Y A0 VDD VDD p L=0.6u W=6u
        M_I$3 Y A0 N$5 GND n L=0.6u W=6u
        M_I$2 N$5 A1 GND GND n L=0.6u W=6u
.ends NAND02_2X

*
* Component pathname : $ADK/parts/nor02_2x
*
.subckt NOR02_2X  A0 A1 Y

        M_I$5 Y A0 GND GND n L=0.6u W=3u
        M_I$4 Y A1 GND GND n L=0.6u W=3u
        M_I$3 Y A1 N$1 VDD p L=0.6u W=7.8u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends NOR02_2X

*
* Component pathname : $ADK/parts/nor03
*
.subckt NOR03  A2 A0 A1 Y

        M_I$213 Y A0 GND GND n L=0.6u W=1.8u
        M_I$211 Y A2 N$211 VDD p L=0.6u W=8.1u
        M_I$5 Y A1 GND GND n L=0.6u W=1.8u
        M_I$4 Y A2 GND GND n L=0.6u W=1.8u
        M_I$3 N$211 A1 N$1 VDD p L=0.6u W=8.1u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=8.1u
.ends NOR03

*
* Component pathname : $ADK/parts/ao21
*
.subckt AO21  A1 A0 B0 Y

        M_I$14 Y N$3 VDD VDD p L=0.6u W=2.7u
        M_I$13 Y N$3 GND GND n L=0.6u W=1.5u
        M_I$12 N$2 A1 GND GND n L=0.6u W=3u
        M_I$11 N$3 A0 N$2 GND n L=0.6u W=3u
        M_I$7 N$3 B0 N$1 VDD p L=0.6u W=3.9u
        M_I$6 N$1 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$1 A0 VDD VDD p L=0.6u W=3.9u
        M_I$4 N$3 B0 GND GND n L=0.6u W=1.5u
.ends AO21

*
* Component pathname : $ADK/parts/mux21
*
.subckt MUX21  S0 A0 A1 Y

        M_I$5 Y S0 N$10 VDD p L=0.6u W=5.4u
        M_I$13 N$6 A1 GND GND n L=0.6u W=3u
        M_I$12 Y S0 N$6 GND n L=0.6u W=3u
        M_I$17 Y N$7 N$5 VDD p L=0.6u W=5.4u
        M_I$16 N$5 A1 VDD VDD p L=0.6u W=5.4u
        M_I$7 N$4 A0 GND GND n L=0.6u W=3u
        M_I$6 Y N$7 N$4 GND n L=0.6u W=3u
        M_I$4 N$10 A0 VDD VDD p L=0.6u W=5.4u
        M_I$3 N$7 S0 GND GND n L=0.6u W=1.5u
        M_I$2 N$7 S0 VDD VDD p L=0.6u W=2.7u
.ends MUX21

*
* Component pathname : /home/max/EECS301/lab3/Areg_S/Areg
*
.subckt AREG  ADDER[0] ADDER[1] ADDER[2] ADDER[3] CONTROL[0] CONTROL[1]
+ A_OUT[0] A_OUT[1] A_OUT[2] A_OUT[3] CLOCK

        X_IX5 NX4 CONTROL[1] CONTROL[0] NAND02_2X
        X_IX11 CONTROL[0] CONTROL[1] NX10 NOR02_2X
        X_IX120 CONTROL[1] NX185 CONTROL[0] NX119 NOR03
        X_IX122 CONTROL[1] A_3 NX119 NX121 AO21
        X_IX181 NX10 CONTROL[1] A_3 ADDER[2] NX180 AOI22
        X_IX175 NX10 CONTROL[1] A_2 ADDER[1] NX174 AOI22
        X_IX169 NX10 CONTROL[1] A_1 ADDER[0] NX168 AOI22
        X_IX186 ADDER[3] NX185 INV02
        X_IX167 CLOCK NOT_CLOCK INV02
        X_IX132 NX4 NX178 NX180 NX131 MUX21
        X_IX142 NX4 NX172 NX174 NX141 MUX21
        X_IX152 NX4 NX164 NX168 NX151 MUX21
        X_REG_AO_3 N$DUMMY_ESC1[4] A_OUT[3] CLOCK A_3 DFF
        X_REG_AO_2 N$DUMMY_ESC1[3] A_OUT[2] CLOCK A_2 DFF
        X_REG_AO_1 N$DUMMY_ESC1[2] A_OUT[1] CLOCK A_1 DFF
        X_REG_A_3 N$DUMMY_ESC1[1] A_3 NOT_CLOCK NX121 DFF
        X_REG_A_2 NX178 A_2 NOT_CLOCK NX131 DFF
        X_REG_A_1 NX172 A_1 NOT_CLOCK NX141 DFF
        X_REG_A_0 NX164 A_0 NOT_CLOCK NX151 DFF
        X_REG_AO_0 N$DUMMY_ESC1[0] A_OUT[0] CLOCK A_0 DFF
.ends AREG

*
* Component pathname : $ADK/parts/oai32
*
.subckt OAI32  A2 B1 A0 A1 B0 Y

        M_I$471 Y A2 N$415 VDD p L=0.6u W=10.8u
        M_I$470 Y A2 N$7 GND n L=0.6u W=4.5u
        M_I$267 N$7 B1 GND GND n L=0.6u W=4.5u
        M_I$265 Y B1 N$414 VDD p L=0.6u W=7.2u
        M_I$5 N$7 B0 GND GND n L=0.6u W=4.5u
        M_I$4 Y A1 N$7 GND n L=0.6u W=4.5u
        M_I$3 Y A0 N$7 GND n L=0.6u W=4.5u
        M_I$12 N$414 B0 VDD VDD p L=0.6u W=7.2u
        M_I$2 N$415 A1 N$9 VDD p L=0.6u W=10.8u
        M_I$1 N$9 A0 VDD VDD p L=0.6u W=10.8u
.ends OAI32

*
* Component pathname : /home/max/EECS301/lab3/Qreg_S/Qreg
*
.subckt QREG  LOAD[0] LOAD[1] LOAD[2] LOAD[3] CONTROL[0] CONTROL[1] Q_OUT[0]
+ Q_OUT[1] Q_OUT[2] Q_OUT[3] Q_OUT[4] A_IN CLOCK

        X_IX5 NX4 CONTROL[1] CONTROL[0] NAND02_2X
        X_IX11 CONTROL[0] CONTROL[1] NX10 NOR02_2X
        X_IX223 NX10 A_IN CONTROL[1] LOAD[3] NX222 AOI22
        X_IX217 NX10 CONTROL[1] Q_4 LOAD[2] NX216 AOI22
        X_IX211 NX10 CONTROL[1] Q_3 LOAD[1] NX210 AOI22
        X_IX203 NX10 CONTROL[1] Q_2 LOAD[0] NX202 AOI22
        X_IX145 NX4 NX220 NX222 NX144 MUX21
        X_IX155 NX4 NX214 NX216 NX154 MUX21
        X_IX165 NX4 NX206 NX210 NX164 MUX21
        X_IX175 NX4 NX199 NX202 NX174 MUX21
        X_IX209 CLOCK NOT_CLOCK INV02
        X_IX198 CONTROL[1] NX197 INV02
        X_IX185 CONTROL[0] NX4 NX197 NX199 NX226 NX184 OAI32
        X_REG_QO_4 N$DUMMY_ESC1[4] Q_OUT[4] CLOCK Q_4 DFF
        X_REG_QO_3 N$DUMMY_ESC1[3] Q_OUT[3] CLOCK Q_3 DFF
        X_REG_QO_2 N$DUMMY_ESC1[2] Q_OUT[2] CLOCK Q_2 DFF
        X_REG_QO_1 N$DUMMY_ESC1[1] Q_OUT[1] CLOCK Q_1 DFF
        X_REG_Q_0 NX226 Q_0 NOT_CLOCK NX184 DFF
        X_REG_Q_4 NX220 Q_4 NOT_CLOCK NX144 DFF
        X_REG_Q_3 NX214 Q_3 NOT_CLOCK NX154 DFF
        X_REG_Q_2 NX206 Q_2 NOT_CLOCK NX164 DFF
        X_REG_Q_1 NX199 Q_1 NOT_CLOCK NX174 DFF
        X_REG_QO_0 N$DUMMY_ESC1[0] Q_OUT[0] CLOCK Q_0 DFF
.ends QREG

*
* Component pathname : $ADK/parts/oai21
*
.subckt OAI21  A0 A1 B0 Y

        M_I$5 N$7 B0 GND GND n L=0.6u W=3u
        M_I$4 Y A1 N$7 GND n L=0.6u W=3u
        M_I$3 Y A0 N$7 GND n L=0.6u W=3u
        M_I$12 Y B0 VDD VDD p L=0.6u W=3.6u
        M_I$2 Y A1 N$9 VDD p L=0.6u W=7.2u
        M_I$1 N$9 A0 VDD VDD p L=0.6u W=7.2u
.ends OAI21

*
* Component pathname : $ADK/parts/nand03
*
.subckt NAND03  A1 Y A0 A2

        M_I$10 Y A2 VDD VDD p L=0.6u W=4.5u
        M_I$9 Y A0 N$4 GND n L=0.6u W=4.5u
        M_I$8 N$5 A2 GND GND n L=0.6u W=4.5u
        M_I$7 N$4 A1 N$5 GND n L=0.6u W=4.5u
        M_I$3 Y A1 VDD VDD p L=0.6u W=4.5u
        M_I$2 Y A0 VDD VDD p L=0.6u W=4.5u
.ends NAND03

*
* Component pathname : $ADK/parts/or02
*
.subckt OR02  A0 A1 Y

        M_I$212 Y N$5 GND GND n L=0.6u W=1.5u
        M_I$211 Y N$5 VDD VDD p L=0.6u W=2.7u
        M_I$5 N$5 A0 GND GND n L=0.6u W=1.5u
        M_I$4 N$5 A1 GND GND n L=0.6u W=1.5u
        M_I$3 N$5 A1 N$1 VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=3.9u
.ends OR02

*
* Component pathname : $ADK/parts/latch
*
.subckt LATCH  Q CLK D

        M_I$222 Q N$17 GND GND n L=0.6u W=1.5u
        M_I$221 Q N$17 VDD VDD p L=0.6u W=2.7u
        M_I$15 N$10 CLK GND GND n L=0.6u W=1.5u
        M_I$13 N$222 N$17 GND GND n L=0.6u W=1.5u
        M_I$12 N$15 N$222 GND GND n L=0.6u W=1.5u
        M_I$11 N$17 N$10 N$15 GND n L=0.6u W=1.5u
        M_I$10 N$13 D GND GND n L=0.6u W=4.5u
        M_I$9 N$17 CLK N$13 GND n L=0.6u W=4.5u
        M_I$6 N$17 CLK N$15 VDD p L=0.6u W=1.5u
        M_I$7 N$222 N$17 VDD VDD p L=0.6u W=2.7u
        M_I$5 N$15 N$222 VDD VDD p L=0.6u W=1.5u
        M_I$4 N$17 N$10 N$11 VDD p L=0.6u W=8.1u
        M_I$3 N$11 D VDD VDD p L=0.6u W=8.1u
        M_I$2 N$10 CLK VDD VDD p L=0.6u W=2.7u
.ends LATCH

*
* Component pathname : $ADK/parts/and03
*
.subckt AND03  A1 Y A0 A2

        M_I$430 Y A VDD VDD p L=0.6u W=2.7u
        M_I$429 Y A GND GND n L=0.6u W=1.5u
        M_I$426 A A2 VDD VDD p L=0.6u W=4.5u
        M_I$425 A A0 N$416 GND n L=0.6u W=4.5u
        M_I$424 N$417 A2 GND GND n L=0.6u W=4.5u
        M_I$423 N$416 A1 N$417 GND n L=0.6u W=4.5u
        M_I$419 A A1 VDD VDD p L=0.6u W=4.5u
        M_I$418 A A0 VDD VDD p L=0.6u W=4.5u
.ends AND03

*
* Component pathname : $ADK/parts/buf02
*
.subckt BUF02  A Y

        M_I$614 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$615 Y N$411 GND GND n L=0.6u W=3u
        M_I$411 N$411 A VDD VDD p L=0.6u W=2.7u
        M_I$412 N$411 A GND GND n L=0.6u W=1.5u
.ends BUF02

*
* Component pathname : $ADK/parts/inv01
*
.subckt INV01  A Y

        M_I$411 Y A VDD VDD p L=0.6u W=2.7u
        M_I$412 Y A GND GND n L=0.6u W=1.5u
.ends INV01

*
* Component pathname : $ADK/parts/latchr
*
.subckt LATCHR  QB R CLK D

        M_I$1954 N$3723 R GND GND n L=0.6u W=3u
        M_I$1953 N$3723 R N$3722 VDD p L=0.6u W=3.6u
        M_I$1244 N$3516 N$3723 VDD VDD p L=0.6u W=1.5u
        M_I$1245 N$3108 N$3723 GND GND n L=0.6u W=1.5u
        M_I$1749 N$3723 N$3929 GND GND n L=0.6u W=3u
        M_I$1240 N$3929 CLK N$3516 VDD p L=0.6u W=1.5u
        M_I$15 N$3100 CLK GND GND n L=0.6u W=1.5u
        M_I$1242 N$3722 N$3929 VDD VDD p L=0.6u W=3.6u
        M_I$1036 QB N$3723 GND GND n L=0.6u W=1.5u
        M_I$10 N$13 D GND GND n L=0.6u W=4.5u
        M_I$9 N$3929 CLK N$13 GND n L=0.6u W=4.5u
        M_I$1035 QB N$3723 VDD VDD p L=0.6u W=2.7u
        M_I$1447 N$3929 N$3100 N$3108 GND n L=0.6u W=1.5u
        M_I$4 N$3929 N$3100 N$11 VDD p L=0.6u W=8.1u
        M_I$3 N$11 D VDD VDD p L=0.6u W=8.1u
        M_I$2 N$3100 CLK VDD VDD p L=0.6u W=2.7u
.ends LATCHR

*
* Component pathname : $ADK/parts/nor02ii
*
.subckt NOR02II  A0 A1 Y

        MP1 N$208 A1 VDD VDD p L=0.6u W=2.7u
        MN1 N$208 A1 GND GND n L=0.6u W=1.5u
        MN4 Y A0 GND GND n L=0.6u W=1.5u
        MN2 Y N$208 GND GND n L=0.6u W=1.5u
        MP4 Y N$208 N$4 VDD p L=0.6u W=3.9u
        MP2 N$4 A0 VDD VDD p L=0.6u W=3.9u
.ends NOR02II

*
* Component pathname : $ADK/parts/buf08
*
.subckt BUF08  A Y

        M_I$1023 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$1022 Y N$411 GND GND n L=0.6u W=3u
        M_I$1021 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$1020 Y N$411 GND GND n L=0.6u W=3u
        M_I$817 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$818 Y N$411 GND GND n L=0.6u W=3u
        M_I$614 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$615 Y N$411 GND GND n L=0.6u W=3u
        M_I$411 N$411 A VDD VDD p L=0.6u W=5.4u
        M_I$412 N$411 A GND GND n L=0.6u W=3u
.ends BUF08

*
* Component pathname : $ADK/parts/inv08
*
.subckt INV08  A Y

        M_I$618 Y A GND GND n L=0.6u W=3u
        M_I$617 Y A VDD VDD p L=0.6u W=5.4u
        M_I$616 Y A GND GND n L=0.6u W=3u
        M_I$619 Y A VDD VDD p L=0.6u W=5.4u
        M_I$412 Y A VDD VDD p L=0.6u W=5.4u
        M_I$413 Y A GND GND n L=0.6u W=3u
        M_I$6 Y A VDD VDD p L=0.6u W=5.4u
        M_I$5 Y A GND GND n L=0.6u W=3u
.ends INV08

*
* Component pathname : $ADK/parts/aoi21
*
.subckt AOI21  A0 A1 B0 Y

        M_I$12 N$8 A1 GND GND n L=0.6u W=3u
        M_I$11 Y A0 N$8 GND n L=0.6u W=3u
        M_I$7 Y B0 N$4 VDD p L=0.6u W=3.9u
        M_I$6 N$4 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$4 A0 VDD VDD p L=0.6u W=3.9u
        M_I$13 Y B0 GND GND n L=0.6u W=1.5u
.ends AOI21

*
* Component pathname : $ADK/parts/nor04
*
.subckt NOR04  A3 A2 A0 A1 Y

        M_I$415 Y A3 GND GND n L=0.6u W=3u
        M_I$416 Y A3 N$418 VDD p L=0.6u W=10.8u
        M_I$213 Y A0 GND GND n L=0.6u W=3u
        M_I$211 N$418 A2 N$211 VDD p L=0.6u W=10.8u
        M_I$5 Y A1 GND GND n L=0.6u W=3u
        M_I$4 Y A2 GND GND n L=0.6u W=3u
        M_I$3 N$211 A1 N$1 VDD p L=0.6u W=10.8u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=10.8u
.ends NOR04

*
* Component pathname : /home/max/EECS301/lab3/Control_S/ControlLogic
*
.subckt CONTROLLOGIC  Q_IN[0] Q_IN[1] Q_SIG[0] Q_SIG[1] A_SIG[0] A_SIG[1]
+ ADDER_SIG M_SIG DONE_SIG START CLOCK

        X_IX129 NX397 NX356 PRES_STATE_0 NX128 NOR03
        X_IX197 PRES_STATE_1 NX440 NX375 NX196 AO21
        X_IX135 COUNT_0 NX411 NX517 NX134 AO21
        X_IX139 NX134 NX128 NX355 NX357 AO21
        X_IX516 NX408 NX517 INV02
        X_IX458 NX517 NX459 INV02
        X_IX439 NX408 NX440 INV02
        X_IX417 NX357 NX416 INV02
        X_IX3 NX414 NX2 INV02
        X_IX429 NX82 NOT_NX82 INV02
        X_IX374 Q_IN[0] NX373 INV02
        X_IX83 NX517 NX72 NX68 NX82 OAI21
        X_IX372 Q_IN[1] NX373 NX375 NX371 OAI21
        X_IX69 NX440 NX68 PRES_STATE_1 PRES_STATE_0 NAND03
        X_IX19 NX414 NX18 NX371 NX416 NAND03
        X_IX415 NX517 NOT_PRES_STATE_0 NX414 OR02
        X_IX53 NEXT_STATE_0 START NX52 OR02
        X_IX147 NEXT_STATE_2 START NX146 OR02
        X_IX31 NEXT_STATE_1 START NX30 OR02
        X_LAT_Q_OUT_1 Q_SIG[1] NX22 NX68 LATCH
        X_LAT_Q_OUT_0 Q_SIG[0] NX22 NOT_NX82 LATCH
        X_LAT_A_OUT_1 A_SIG[1] NX22 NOT_PRES_STATE_0 LATCH
        X_LAT_A_OUT_0 A_SIG[0] NX444 NX196 LATCH
        X_LAT_DONE DONE_SIG NX444 NX355 LATCH
        X_LAT_M_OUT M_SIG NX444 PRES_STATE_0 LATCH
        X_LAT_COUNT_0 COUNT_0 NX446 NX94 LATCH
        X_LAT_NEXT_STATE_0 NEXT_STATE_0 NX444 NX44 LATCH
        X_LAT_COUNT_2 COUNT_2 NX446 NX356 LATCH
        X_LAT_NEXT_STATE_2 NEXT_STATE_2 NX444 NX357 LATCH
        X_LAT_NEXT_STATE_1 NEXT_STATE_1 NX444 NX18 LATCH
        X_LAT_ADDER ADDER_SIG NX2 PRES_STATE_1 LATCH
        X_IX111 NX406 NX440 NX110 NOR02_2X
        X_IX95 COUNT_0 NX440 NX94 NOR02_2X
        X_IX157 NOT_PRES_STATE_0 NX355 NX517 PRES_STATE_1 AND03
        X_IX456 NX400 NX457 BUF02
        X_LAT_COUNT_1__U3 NX5 NX411 BUF02
        X_LAT_COUNT_1__U2 NX5 COUNT_1 INV01
        X_LAT_COUNT_1__U1 NX5 GND NX446 NX448 LATCHR
        X_IX401 COUNT_0 NX411 NX400 NOR02II
        X_IX447 NX110 NX448 BUF08
        X_IX445 NOT_NX82 NX446 INV08
        X_IX407 COUNT_1 COUNT_0 NX457 NX406 AOI21
        X_REG_PRES_STATE_2 NX408 N$DUMMY_ESC1[0] CLOCK NX146 DFF
        X_REG_PRES_STATE_1 NX397 PRES_STATE_1 CLOCK NX30 DFF
        X_REG_PRES_STATE_0 NOT_PRES_STATE_0 PRES_STATE_0 CLOCK NX52 DFF
        X_IX45 NX394 PRES_STATE_0 PRES_STATE_1 NX517 NX44 NOR04
        X_IX395 NX394 Q_IN[1] Q_IN[0] XNOR2
        X_IX384 NX383 COUNT_2 NX457 XNOR2
        X_IX443 NX444 NX397 NX440 NAND02_2X
        X_IX23 NX22 NX397 NX440 NAND02_2X
        X_IX73 NX72 NOT_PRES_STATE_0 PRES_STATE_1 NAND02_2X
        X_IX123 NX356 NX383 NX459 NAND02_2X
        X_IX376 PRES_STATE_0 PRES_STATE_1 NX517 NX375 NOR03
.ends CONTROLLOGIC

*
* MAIN CELL: Component pathname : /home/max/EECS301/lab3/TopModel
*
        X_ADDSUB1 N$1[0] N$1[1] N$1[2] N$1[3] OUT[4] OUT[5] OUT[6] OUT[7]
+ N$2[0] N$2[1] N$2[2] N$2[3] CLK ADDCONTROL ADDSUB
        X_MREG1 MIN[0] MIN[1] MIN[2] MIN[3] N$1[0] N$1[1] N$1[2] N$1[3]
+ CLK N$62 MREG
        X_AREG1 N$2[0] N$2[1] N$2[2] N$2[3] ACONTROL[0] ACONTROL[1] OUT[4]
+ OUT[5] OUT[6] OUT[7] CLK AREG
        X_QREG1 QIN[0] QIN[1] QIN[2] QIN[3] QCONTROL[0] QCONTROL[1] Q[0]
+ OUT[0] OUT[1] OUT[2] OUT[3] OUT[4] CLK QREG
        X_CONTROLLOGIC1 Q[0] OUT[0] QCONTROL[0] QCONTROL[1] ACONTROL[0]
+ ACONTROL[1] ADDCONTROL N$62 DONE START CLK CONTROLLOGIC
*
.end
