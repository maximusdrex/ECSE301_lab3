*
* .CONNECT statements
*
.CONNECT GND 0


* ELDO netlist generated with ICnet by 'max' on Mon Mar 21 2022 at 13:20:18

*
* Globals.
*
.global VDD GND

*
* Component pathname : $ADK/parts/latch
*
.subckt LATCH  Q CLK D

        M_I$222 Q N$17 GND GND n L=0.6u W=1.5u
        M_I$221 Q N$17 VDD VDD p L=0.6u W=2.7u
        M_I$15 N$10 CLK GND GND n L=0.6u W=1.5u
        M_I$13 N$222 N$17 GND GND n L=0.6u W=1.5u
        M_I$12 N$15 N$222 GND GND n L=0.6u W=1.5u
        M_I$11 N$17 N$10 N$15 GND n L=0.6u W=1.5u
        M_I$10 N$13 D GND GND n L=0.6u W=4.5u
        M_I$9 N$17 CLK N$13 GND n L=0.6u W=4.5u
        M_I$6 N$17 CLK N$15 VDD p L=0.6u W=1.5u
        M_I$7 N$222 N$17 VDD VDD p L=0.6u W=2.7u
        M_I$5 N$15 N$222 VDD VDD p L=0.6u W=1.5u
        M_I$4 N$17 N$10 N$11 VDD p L=0.6u W=8.1u
        M_I$3 N$11 D VDD VDD p L=0.6u W=8.1u
        M_I$2 N$10 CLK VDD VDD p L=0.6u W=2.7u
.ends LATCH

*
* Component pathname : $ADK/parts/buf02
*
.subckt BUF02  A Y

        M_I$614 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$615 Y N$411 GND GND n L=0.6u W=3u
        M_I$411 N$411 A VDD VDD p L=0.6u W=2.7u
        M_I$412 N$411 A GND GND n L=0.6u W=1.5u
.ends BUF02

*
* Component pathname : $ADK/parts/inv02
*
.subckt INV02  A Y

        M_I$6 Y A VDD VDD p L=0.6u W=5.4u
        M_I$5 Y A GND GND n L=0.6u W=3u
.ends INV02

*
* Component pathname : $ADK/parts/nand02_2x
*
.subckt NAND02_2X  Y A0 A1

        M_I$9 Y A1 VDD VDD p L=0.6u W=6u
        M_I$8 Y A0 VDD VDD p L=0.6u W=6u
        M_I$3 Y A0 N$5 GND n L=0.6u W=6u
        M_I$2 N$5 A1 GND GND n L=0.6u W=6u
.ends NAND02_2X

*
* Component pathname : $ADK/parts/nor02_2x
*
.subckt NOR02_2X  A0 A1 Y

        M_I$5 Y A0 GND GND n L=0.6u W=3u
        M_I$4 Y A1 GND GND n L=0.6u W=3u
        M_I$3 Y A1 N$1 VDD p L=0.6u W=7.8u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends NOR02_2X

*
* Component pathname : $ADK/parts/xnor2
*
.subckt XNOR2  Y A0 A1

        M_I$218 N$213 A1 GND GND n L=0.6u W=3u
        M_I$217 N$212 A0 N$213 GND n L=0.6u W=3u
        M_I$9 N$212 A1 VDD VDD p L=0.6u W=3.9u
        M_I$8 N$212 A0 VDD VDD p L=0.6u W=3.9u
        M_I$7 N$3 N$212 GND GND n L=0.6u W=3u
        M_I$6 Y A1 N$3 GND n L=0.6u W=3u
        M_I$5 Y A0 N$3 GND n L=0.6u W=3u
        M_I$4 Y A1 N$1 VDD p L=0.6u W=7.8u
        M_I$3 Y N$212 VDD VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends XNOR2

*
* Component pathname : $ADK/parts/nor03
*
.subckt NOR03  A2 A0 A1 Y

        M_I$213 Y A0 GND GND n L=0.6u W=1.8u
        M_I$211 Y A2 N$211 VDD p L=0.6u W=8.1u
        M_I$5 Y A1 GND GND n L=0.6u W=1.8u
        M_I$4 Y A2 GND GND n L=0.6u W=1.8u
        M_I$3 N$211 A1 N$1 VDD p L=0.6u W=8.1u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=8.1u
.ends NOR03

*
* Component pathname : $ADK/parts/ao21
*
.subckt AO21  A1 A0 B0 Y

        M_I$14 Y N$3 VDD VDD p L=0.6u W=2.7u
        M_I$13 Y N$3 GND GND n L=0.6u W=1.5u
        M_I$12 N$2 A1 GND GND n L=0.6u W=3u
        M_I$11 N$3 A0 N$2 GND n L=0.6u W=3u
        M_I$7 N$3 B0 N$1 VDD p L=0.6u W=3.9u
        M_I$6 N$1 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$1 A0 VDD VDD p L=0.6u W=3.9u
        M_I$4 N$3 B0 GND GND n L=0.6u W=1.5u
.ends AO21

*
* Component pathname : $ADK/parts/dff
*
.subckt DFF  QB Q CLK D

        M_I$441 N$847 BCLK- N$851 GND n L=0.6u W=4.5u
        M_I$440 N$849 N$847 VDD VDD p L=0.6u W=1.5u
        M_I$439 N$847 BCLK- N$848 VDD p L=0.6u W=1.5u
        M_I$438 N$848 N$849 VDD VDD p L=0.6u W=1.5u
        M_I$437 N$847 BCLK N$845 VDD p L=0.6u W=8.1u
        M_I$436 N$845 D VDD VDD p L=0.6u W=8.1u
        M_I$452 BCLK BCLK- GND GND n L=0.6u W=3u
        M_I$673 Q QB GND GND n L=0.6u W=3u
        M_I$672 Q QB VDD VDD p L=0.6u W=5.4u
        M_I$669 QB N$1074 GND GND n L=0.6u W=3u
        M_I$675 QB N$1074 VDD VDD p L=0.6u W=5.4u
        M_I$668 N$1071 N$1074 GND GND n L=0.6u W=1.5u
        M_I$667 N$1073 N$1071 GND GND n L=0.6u W=1.5u
        M_I$666 N$1074 BCLK- N$1073 GND n L=0.6u W=1.5u
        M_I$665 N$1072 N$847 GND GND n L=0.6u W=4.5u
        M_I$664 N$1074 BCLK N$1072 GND n L=0.6u W=4.5u
        M_I$663 N$1071 N$1074 VDD VDD p L=0.6u W=1.5u
        M_I$662 N$1074 BCLK N$1070 VDD p L=0.6u W=1.5u
        M_I$661 N$1070 N$1071 VDD VDD p L=0.6u W=1.5u
        M_I$660 N$1074 BCLK- N$1069 VDD p L=0.6u W=8.1u
        M_I$659 N$1069 N$847 VDD VDD p L=0.6u W=8.1u
        M_I$449 BCLK- CLK GND GND n L=0.6u W=3u
        M_I$448 BCLK- CLK VDD VDD p L=0.6u W=5.4u
        M_I$453 BCLK BCLK- VDD VDD p L=0.6u W=5.4u
        M_I$445 N$849 N$847 GND GND n L=0.6u W=1.5u
        M_I$444 N$852 N$849 GND GND n L=0.6u W=1.5u
        M_I$443 N$847 BCLK N$852 GND n L=0.6u W=1.5u
        M_I$442 N$851 D GND GND n L=0.6u W=4.5u
.ends DFF

*
* Component pathname : $ADK/parts/and02
*
.subckt AND02  Y A0 A1

        M_I$674 Y N$5 VDD VDD p L=0.6u W=2.7u
        M_I$675 Y N$5 GND GND n L=0.6u W=1.5u
        M_I$472 N$5 A1 VDD VDD p L=0.6u W=3.6u
        M_I$471 N$5 A0 VDD VDD p L=0.6u W=3.6u
        M_I$4 N$5 A0 N$7 GND n L=0.6u W=3u
        M_I$5 N$7 A1 GND GND n L=0.6u W=3u
.ends AND02

*
* Component pathname : $ADK/parts/oai21
*
.subckt OAI21  A0 A1 B0 Y

        M_I$5 N$7 B0 GND GND n L=0.6u W=3u
        M_I$4 Y A1 N$7 GND n L=0.6u W=3u
        M_I$3 Y A0 N$7 GND n L=0.6u W=3u
        M_I$12 Y B0 VDD VDD p L=0.6u W=3.6u
        M_I$2 Y A1 N$9 VDD p L=0.6u W=7.2u
        M_I$1 N$9 A0 VDD VDD p L=0.6u W=7.2u
.ends OAI21

*
* Component pathname : $ADK/parts/inv01
*
.subckt INV01  A Y

        M_I$411 Y A VDD VDD p L=0.6u W=2.7u
        M_I$412 Y A GND GND n L=0.6u W=1.5u
.ends INV01

*
* Component pathname : $ADK/parts/latchr
*
.subckt LATCHR  QB R CLK D

        M_I$1954 N$3723 R GND GND n L=0.6u W=3u
        M_I$1953 N$3723 R N$3722 VDD p L=0.6u W=3.6u
        M_I$1244 N$3516 N$3723 VDD VDD p L=0.6u W=1.5u
        M_I$1245 N$3108 N$3723 GND GND n L=0.6u W=1.5u
        M_I$1749 N$3723 N$3929 GND GND n L=0.6u W=3u
        M_I$1240 N$3929 CLK N$3516 VDD p L=0.6u W=1.5u
        M_I$15 N$3100 CLK GND GND n L=0.6u W=1.5u
        M_I$1242 N$3722 N$3929 VDD VDD p L=0.6u W=3.6u
        M_I$1036 QB N$3723 GND GND n L=0.6u W=1.5u
        M_I$10 N$13 D GND GND n L=0.6u W=4.5u
        M_I$9 N$3929 CLK N$13 GND n L=0.6u W=4.5u
        M_I$1035 QB N$3723 VDD VDD p L=0.6u W=2.7u
        M_I$1447 N$3929 N$3100 N$3108 GND n L=0.6u W=1.5u
        M_I$4 N$3929 N$3100 N$11 VDD p L=0.6u W=8.1u
        M_I$3 N$11 D VDD VDD p L=0.6u W=8.1u
        M_I$2 N$3100 CLK VDD VDD p L=0.6u W=2.7u
.ends LATCHR

*
* Component pathname : $ADK/parts/or03
*
.subckt OR03  A2 A0 A1 Y

        M_I$416 Y N$214 GND GND n L=0.6u W=1.5u
        M_I$415 Y N$214 VDD VDD p L=0.6u W=2.7u
        M_I$213 N$214 A0 GND GND n L=0.6u W=1.8u
        M_I$211 N$214 A2 N$211 VDD p L=0.6u W=8.1u
        M_I$5 N$214 A1 GND GND n L=0.6u W=1.8u
        M_I$4 N$214 A2 GND GND n L=0.6u W=1.8u
        M_I$3 N$211 A1 N$1 VDD p L=0.6u W=8.1u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=8.1u
.ends OR03

*
* Component pathname : $ADK/parts/buf08
*
.subckt BUF08  A Y

        M_I$1023 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$1022 Y N$411 GND GND n L=0.6u W=3u
        M_I$1021 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$1020 Y N$411 GND GND n L=0.6u W=3u
        M_I$817 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$818 Y N$411 GND GND n L=0.6u W=3u
        M_I$614 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$615 Y N$411 GND GND n L=0.6u W=3u
        M_I$411 N$411 A VDD VDD p L=0.6u W=5.4u
        M_I$412 N$411 A GND GND n L=0.6u W=3u
.ends BUF08

*
* Component pathname : $ADK/parts/inv08
*
.subckt INV08  A Y

        M_I$618 Y A GND GND n L=0.6u W=3u
        M_I$617 Y A VDD VDD p L=0.6u W=5.4u
        M_I$616 Y A GND GND n L=0.6u W=3u
        M_I$619 Y A VDD VDD p L=0.6u W=5.4u
        M_I$412 Y A VDD VDD p L=0.6u W=5.4u
        M_I$413 Y A GND GND n L=0.6u W=3u
        M_I$6 Y A VDD VDD p L=0.6u W=5.4u
        M_I$5 Y A GND GND n L=0.6u W=3u
.ends INV08

*
* Component pathname : $ADK/parts/nor03_2x
*
.subckt NOR03_2X  A1 A0 A2 Y

        M_I$12 Y A0 GND GND n L=0.6u W=3.3u
        M_I$10 Y A2 N$3 VDD p L=0.6u W=12u
        M_I$5 Y A1 GND GND n L=0.6u W=3.3u
        M_I$4 Y A2 GND GND n L=0.6u W=3.3u
        M_I$3 N$3 A1 N$1 VDD p L=0.6u W=12u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=12u
.ends NOR03_2X

*
* Component pathname : $ADK/parts/nor04
*
.subckt NOR04  A3 A2 A0 A1 Y

        M_I$415 Y A3 GND GND n L=0.6u W=3u
        M_I$416 Y A3 N$418 VDD p L=0.6u W=10.8u
        M_I$213 Y A0 GND GND n L=0.6u W=3u
        M_I$211 N$418 A2 N$211 VDD p L=0.6u W=10.8u
        M_I$5 Y A1 GND GND n L=0.6u W=3u
        M_I$4 Y A2 GND GND n L=0.6u W=3u
        M_I$3 N$211 A1 N$1 VDD p L=0.6u W=10.8u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=10.8u
.ends NOR04

*
* Component pathname : $ADK/parts/or02
*
.subckt OR02  A0 A1 Y

        M_I$212 Y N$5 GND GND n L=0.6u W=1.5u
        M_I$211 Y N$5 VDD VDD p L=0.6u W=2.7u
        M_I$5 N$5 A0 GND GND n L=0.6u W=1.5u
        M_I$4 N$5 A1 GND GND n L=0.6u W=1.5u
        M_I$3 N$5 A1 N$1 VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=3.9u
.ends OR02

*
* Component pathname : $ADK/parts/nor02ii
*
.subckt NOR02II  A0 A1 Y

        MP1 N$208 A1 VDD VDD p L=0.6u W=2.7u
        MN1 N$208 A1 GND GND n L=0.6u W=1.5u
        MN4 Y A0 GND GND n L=0.6u W=1.5u
        MN2 Y N$208 GND GND n L=0.6u W=1.5u
        MP4 Y N$208 N$4 VDD p L=0.6u W=3.9u
        MP2 N$4 A0 VDD VDD p L=0.6u W=3.9u
.ends NOR02II

*
* Component pathname : $ADK/parts/ao22
*
.subckt AO22  A1 A0 B0 Y B1

        M_I$16 Y N$215 VDD VDD p L=0.6u W=2.7u
        M_I$18 Y N$215 GND GND n L=0.6u W=1.5u
        M_I$14 N$215 B0 N$2 GND n L=0.6u W=3u
        M_I$13 N$215 B1 N$6 VDD p L=0.6u W=3.9u
        M_I$12 N$1 A1 GND GND n L=0.6u W=3u
        M_I$11 N$215 A0 N$1 GND n L=0.6u W=3u
        M_I$7 N$215 B0 N$6 VDD p L=0.6u W=3.9u
        M_I$6 N$6 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$6 A0 VDD VDD p L=0.6u W=3.9u
        M_I$4 N$2 B1 GND GND n L=0.6u W=3u
.ends AO22

*
* Component pathname : $ADK/parts/mux21_ni
*
.subckt MUX21_NI  S0 A0 A1 Y

        M_I$18 Y N$11 GND GND n L=0.6u W=1.5u
        M_I$17 Y N$11 VDD VDD p L=0.6u W=2.7u
        M_I$16 N$11 S0 N$7 VDD p L=0.6u W=5.4u
        M_I$11 N$3 A1 GND GND n L=0.6u W=3u
        M_I$10 N$11 S0 N$3 GND n L=0.6u W=3u
        M_I$9 N$11 N$4 N$2 VDD p L=0.6u W=5.4u
        M_I$8 N$2 A1 VDD VDD p L=0.6u W=5.4u
        M_I$7 N$1 A0 GND GND n L=0.6u W=3u
        M_I$6 N$11 N$4 N$1 GND n L=0.6u W=3u
        M_I$4 N$7 A0 VDD VDD p L=0.6u W=5.4u
        M_I$3 N$4 S0 GND GND n L=0.6u W=1.5u
        M_I$2 N$4 S0 VDD VDD p L=0.6u W=2.7u
.ends MUX21_NI

*
* Component pathname : $ADK/parts/ao32
*
.subckt AO32  Y A0 A1 A2 B0 B1

        M_I$222 Y N$214 GND GND n L=0.6u W=1.5u
        M_I$221 Y N$214 VDD VDD p L=0.6u W=2.7u
        M_I$12 N$6 B1 GND GND n L=0.6u W=3u
        M_I$11 N$214 B0 N$6 GND n L=0.6u W=3u
        M_I$10 N$5 A2 GND GND n L=0.6u W=4.5u
        M_I$9 N$4 A1 N$5 GND n L=0.6u W=4.5u
        M_I$8 N$214 A0 N$4 GND n L=0.6u W=4.5u
        M_I$6 N$214 B0 N$11 VDD p L=0.6u W=3.9u
        M_I$5 N$214 B1 N$11 VDD p L=0.6u W=3.9u
        M_I$4 N$11 A0 VDD VDD p L=0.6u W=3.9u
        M_I$3 N$11 A1 VDD VDD p L=0.6u W=3.9u
        M_I$2 N$11 A2 VDD VDD p L=0.6u W=3.9u
.ends AO32

*
* Component pathname : $ADK/parts/xor2
*
.subckt XOR2  Y A0 A1

        M_I$421 Y N$4 GND GND n L=0.6u W=1.5u
        M_I$420 Y N$4 VDD VDD p L=0.6u W=2.7u
        M_I$218 N$213 A1 GND GND n L=0.6u W=3u
        M_I$217 N$212 A0 N$213 GND n L=0.6u W=3u
        M_I$9 N$212 A1 VDD VDD p L=0.6u W=3.9u
        M_I$8 N$212 A0 VDD VDD p L=0.6u W=3.9u
        M_I$7 N$3 N$212 GND GND n L=0.6u W=3u
        M_I$6 N$4 A1 N$3 GND n L=0.6u W=3u
        M_I$5 N$4 A0 N$3 GND n L=0.6u W=3u
        M_I$4 N$4 A1 N$1 VDD p L=0.6u W=7.8u
        M_I$3 N$4 N$212 VDD VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends XOR2

*
* Component pathname : $ADK/parts/aoi22
*
.subckt AOI22  B1 A0 A1 B0 Y

        M_I$425 Y B0 N$9 GND n L=0.6u W=3u
        M_I$426 Y B1 N$4 VDD p L=0.6u W=3.9u
        M_I$12 N$8 A1 GND GND n L=0.6u W=3u
        M_I$11 Y A0 N$8 GND n L=0.6u W=3u
        M_I$7 Y B0 N$4 VDD p L=0.6u W=3.9u
        M_I$6 N$4 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$4 A0 VDD VDD p L=0.6u W=3.9u
        M_I$13 N$9 B1 GND GND n L=0.6u W=3u
.ends AOI22

*
* MAIN CELL: Component pathname : /home/max/301/ECSE301_lab3/TopModel_S/TopModel
*
        X_CONTROL_LAT_COUNT_1 CONTROL_COUNT_1 CONTROL_NX14 CONTROL_NX80 LATCH
        X_CONTROL_LAT_COUNT_2 CONTROL_COUNT_2 CONTROL_NX14 CONTROL_NX108 LATCH
        X_CONTROL_LAT_ADDER_SIG ADD_SIG CONTROL_NX646 CONTROL_PRES_STATE_2 LATCH
        X_CONTROL_LAT_NEXT_STATE_3 CONTROL_NEXT_STATE_3 CONTROL_NX646 CONTROL_NX62 LATCH
        X_CONTROL_LAT_M_SIG M_SIG CONTROL_NX648 CONTROL_PRES_STATE_4 LATCH
        X_CONTROL_LAT_Q_SIG_0 Q_CON_0 CONTROL_NX648 CONTROL_NX10 LATCH
        X_CONTROL_LAT_NEXT_STATE_2 CONTROL_NEXT_STATE_2 CONTROL_NX646 CONTROL_NX190 LATCH
        X_CONTROL_LAT_NEXT_STATE_0 CONTROL_NEXT_STATE_0 CONTROL_NX646 CONTROL_NX168 LATCH
        X_CONTROL_IX645 CONTROL_NX36 CONTROL_NX646 BUF02
        X_CONTROL_IX647 CONTROL_NX36 CONTROL_NX648 BUF02
        X_IX371 A_CON_1 NX372 BUF02
        X_IX373 A_CON_1 NX374 BUF02
        X_CONTROL_LAT_COUNT_0__U3 CONTROL_NX5 CONTROL_NX622 BUF02
        X_CONTROL_IX660 CONTROL_NX609 CONTROL_NX661 BUF02
        X_CONTROL_IX29 CONTROL_NX592 CONTROL_NX28 INV02
        X_CONTROL_IX617 CLOCK CONTROL_NX616 INV02
        X_CONTROL_IX37 CONTROL_NX36 CONTROL_NX590 CONTROL_NX625 NAND02_2X
        X_CONTROL_IX151 START CONTROL_NX598 CONTROL_NX150 NOR02_2X
        X_CONTROL_IX11 CONTROL_PRES_STATE_4 CONTROL_PRES_STATE_3 CONTROL_NX10 NOR02_2X
        X_CONTROL_IX608 CONTROL_NX607 CONTROL_COUNT_2 CONTROL_NX661 XNOR2
        X_CONTROL_IX593 CONTROL_PRES_STATE_0 CONTROL_PRES_STATE_4 CONTROL_PRES_STATE_5
+ CONTROL_NX592 NOR03
        X_CONTROL_IX191 Q_OUT_0 CONTROL_NX569 CONTROL_NX630 CONTROL_NX190 NOR03
        X_CONTROL_IX131 CONTROL_PRES_STATE_5 START CONTROL_NX126 CONTROL_NX130 AO21
        X_CONTROL_IX591 CONTROL_NX24 CONTROL_NX592 CONTROL_NX616 CONTROL_NX590 AO21
        X_CONTROL_IX61 CONTROL_NX581 CONTROL_PRES_STATE_0 CONTROL_PRES_STATE_1
+ CONTROL_NX60 AO21
        X_CONTROL_IX105 CONTROL_COUNT_0 CONTROL_COUNT_1 CONTROL_NX661 CONTROL_NX556 AO21
        X_CONTROL_IX169 CONTROL_NX656 CONTROL_PRES_STATE_3 CONTROL_PRES_STATE_4
+ CONTROL_NX168 AO21
        X_CONTROL_REG_PRES_STATE_5 CONTROL_NX598 CONTROL_PRES_STATE_5 CLOCK
+ CONTROL_NX140 DFF
        X_CONTROL_REG_PRES_STATE_4 CONTROL_NOT_PRES_STATE_4 CONTROL_PRES_STATE_4
+ CLOCK CONTROL_NX158 DFF
        X_CONTROL_REG_PRES_STATE_3 CONTROL_NX574 CONTROL_PRES_STATE_3 CLOCK
+ CONTROL_NX72 DFF
        X_CONTROL_REG_PRES_STATE_0 CONTROL_NX569 CONTROL_PRES_STATE_0 CLOCK
+ CONTROL_NX178 DFF
        X_CONTROL_IX81 CONTROL_NX80 CONTROL_PRES_STATE_3 CONTROL_NX556 AND02
        X_CONTROL_IX109 CONTROL_NX574 CONTROL_NX607 CONTROL_NOT_PRES_STATE_4
+ CONTROL_NX108 OAI21
        X_CONTROL_IX626 CONTROL_PRES_STATE_4 CONTROL_PRES_STATE_3 CLOCK
+ CONTROL_NX625 OAI21
        X_CONTROL_LAT_COUNT_0__U2 CONTROL_NX5 CONTROL_COUNT_0 INV01
        X_CONTROL_LAT_COUNT_0__U1 CONTROL_NX5 GND CONTROL_NX14 CONTROL_NX650 LATCHR
        X_CONTROL_IX629 CONTROL_COUNT_1 CONTROL_COUNT_2 CONTROL_NX622 CONTROL_NX656 OR03
        X_CONTROL_IX649 CONTROL_NX90 CONTROL_NX650 BUF08
        X_CONTROL_IX15 CONTROL_NX625 CONTROL_NX14 INV08
        X_CONTROL_IX25 CONTROL_PRES_STATE_4 CONTROL_PRES_STATE_1 CONTROL_PRES_STATE_2
+ CONTROL_NX24 NOR03_2X
        X_CONTROL_IX127 CONTROL_COUNT_1 CONTROL_NX622 CONTROL_NX574 CONTROL_COUNT_2
+ CONTROL_NX126 NOR04
        X_CONTROL_IX159 CONTROL_NEXT_STATE_4 START CONTROL_NX158 OR02
        X_CONTROL_IX63 CONTROL_NX60 CONTROL_PRES_STATE_2 CONTROL_NX62 OR02
        X_CONTROL_IX141 START CONTROL_NEXT_STATE_5 CONTROL_NX140 NOR02II
        X_CONTROL_IX47 START CONTROL_NEXT_STATE_1 CONTROL_NX46 NOR02II
        X_CONTROL_IX91 CONTROL_NX574 CONTROL_NX622 CONTROL_NX90 NOR02II
        X_CONTROL_IX610 CONTROL_COUNT_1 CONTROL_NX622 CONTROL_NX609 NOR02II
        X_CONTROL_IX73 START CONTROL_NEXT_STATE_3 CONTROL_NX72 NOR02II
        X_CONTROL_IX201 START CONTROL_NEXT_STATE_2 CONTROL_NX200 NOR02II
        X_CONTROL_IX179 START CONTROL_NEXT_STATE_0 CONTROL_NX178 NOR02II
        X_CONTROL_LAT_NEXT_STATE_5 CONTROL_NEXT_STATE_5 CONTROL_NX646 CONTROL_NX130 LATCH
        X_CONTROL_LAT_NEXT_STATE_1 CONTROL_NEXT_STATE_1 CONTROL_NX646 CONTROL_NX4 LATCH
        X_CONTROL_LAT_NEXT_STATE_4 CONTROL_NEXT_STATE_4 CONTROL_NX646 CONTROL_NX150 LATCH
        X_CONTROL_LAT_A_SIG_0 A_CON_0 CONTROL_NX648 CONTROL_NX28 LATCH
        X_CONTROL_LAT_Q_SIG_1 Q_CON_1 CONTROL_NX648 CONTROL_NOT_PRES_STATE_4 LATCH
        X_CONTROL_LAT_DONE_SIG DONE CONTROL_NX648 CONTROL_PRES_STATE_5 LATCH
        X_CONTROL_LAT_A_SIG_1 A_CON_1 CONTROL_NX648 CONTROL_NX24 LATCH
        X_IX357 CLOCK NOT_CLOCK INV02
        X_IX310 NX309 NX311 NX332 XNOR2
        X_IX87 NX86 NX341 NX84 XNOR2
        X_IX83 NX82 ADD_SIG M_OUT_2 XNOR2
        X_IX61 NX60 ADD_SIG M_OUT_1 XNOR2
        X_CONTROL_IX582 CONTROL_NX581 MULT_OUT[0] Q_OUT_0 XNOR2
        X_IX352 NX351 M_OUT_0 MULT_OUT[4] XNOR2
        X_IX63 NX62 NX60 MULT_OUT[5] XNOR2
        X_IX85 NX84 NX82 MULT_OUT[6] XNOR2
        X_IX333 NX332 MULT_OUT[7] NX334 XNOR2
        X_IX45 NX374 NX351 A_CON_0 NX44 NOR03
        X_IX67 NX374 NX347 A_CON_0 NX66 NOR03
        X_IX192 NX372 A_CON_0 NX309 NX191 NOR03
        X_CONTROL_IX5 CONTROL_NX587 CONTROL_NX569 MULT_OUT[0] CONTROL_NX4 NOR03
        X_IX145 MULT_OUT[5] NX372 NX44 NX144 AO21
        X_IX135 MULT_OUT[6] NX372 NX66 NX134 AO21
        X_IX194 NX372 MULT_OUT[7] NX191 NX193 AO21
        X_IX187 MULT_OUT[1] Q_CON_1 Q_IN[0] NX186 NX10 AO22
        X_IX204 NX24 MULT_OUT[6] NX124 NX203 MUX21_NI
        X_IX274 NX273 Q_CON_1 MULT_OUT[0] NX362 Q_OUT_0 NX364 AO32
        X_CONTROL_REG_PRES_STATE_1 N$DUMMY_ESC1[14] CONTROL_PRES_STATE_1
+ CLOCK CONTROL_NX46 DFF
        X_CONTROL_REG_PRES_STATE_2 N$DUMMY_ESC1[13] CONTROL_PRES_STATE_2
+ CLOCK CONTROL_NX200 DFF
        X_M_REG_M_OUT_3 N$DUMMY_ESC1[12] M_OUT_3 CLOCK NX183 DFF
        X_M_REG_M_OUT_1 N$DUMMY_ESC1[11] M_OUT_1 CLOCK NX163 DFF
        X_M_REG_M_OUT_0 N$DUMMY_ESC1[10] M_OUT_0 CLOCK NX153 DFF
        X_M_REG_M_OUT_2 N$DUMMY_ESC1[9] M_OUT_2 CLOCK NX173 DFF
        X_A_REG_A_OUT_3 N$DUMMY_ESC1[8] MULT_OUT[7] CLOCK NX193 DFF
        X_A_REG_A_OUT_2 N$DUMMY_ESC1[7] MULT_OUT[6] CLOCK NX203 DFF
        X_A_REG_A_OUT_1 N$DUMMY_ESC1[6] MULT_OUT[5] CLOCK NX213 DFF
        X_A_REG_A_OUT_0 N$DUMMY_ESC1[5] MULT_OUT[4] CLOCK NX223 DFF
        X_Q_REG_Q_OUT_4 N$DUMMY_ESC1[4] MULT_OUT[3] NOT_CLOCK NX233 DFF
        X_Q_REG_Q_OUT_3 N$DUMMY_ESC1[3] MULT_OUT[2] NOT_CLOCK NX243 DFF
        X_Q_REG_Q_OUT_2 N$DUMMY_ESC1[2] MULT_OUT[1] NOT_CLOCK NX253 DFF
        X_Q_REG_Q_OUT_1 N$DUMMY_ESC1[1] MULT_OUT[0] NOT_CLOCK NX263 DFF
        X_Q_REG_Q_OUT_0 N$DUMMY_ESC1[0] Q_OUT_0 NOT_CLOCK NX273 DFF
        X_IX363 Q_CON_0 NX362 INV02
        X_CONTROL_IX588 Q_OUT_0 CONTROL_NX587 INV02
        X_IX365 NX4 NX364 INV02
        X_IX329 NX60 NX328 INV02
        X_IX75 NX341 NX74 INV02
        X_IX314 NX82 NX313 INV02
        X_CONTROL_IX631 MULT_OUT[0] CONTROL_NX630 INV02
        X_IX5 NX4 Q_CON_1 Q_CON_0 NAND02_2X
        X_IX25 NX24 NX372 A_CON_0 NAND02_2X
        X_IX11 Q_CON_0 Q_CON_1 NX10 NOR02_2X
        X_IX43 A_CON_0 NX372 NX42 NOR02_2X
        X_IX335 NX334 ADD_SIG M_OUT_3 XOR2
        X_IX342 MULT_OUT[5] NX52 NX62 NX328 NX341 AOI22
        X_IX312 NX84 NX313 MULT_OUT[6] NX74 NX311 AOI22
        X_IX348 NX347 NX52 NX62 XNOR2
        X_IX177 MULT_OUT[2] Q_CON_1 Q_IN[1] NX176 NX10 AO22
        X_IX167 MULT_OUT[3] Q_CON_1 Q_IN[2] NX166 NX10 AO22
        X_IX155 MULT_OUT[4] Q_CON_1 Q_IN[3] NX154 NX10 AO22
        X_IX125 MULT_OUT[7] NX372 NX86 NX124 NX42 AO22
        X_IX154 M_SIG M_OUT_0 M_IN[0] NX153 MUX21_NI
        X_IX164 M_SIG M_OUT_1 M_IN[1] NX163 MUX21_NI
        X_IX174 M_SIG M_OUT_2 M_IN[2] NX173 MUX21_NI
        X_IX184 M_SIG M_OUT_3 M_IN[3] NX183 MUX21_NI
        X_IX264 NX4 MULT_OUT[0] NX186 NX263 MUX21_NI
        X_IX254 NX4 MULT_OUT[1] NX176 NX253 MUX21_NI
        X_IX244 NX4 MULT_OUT[2] NX166 NX243 MUX21_NI
        X_IX234 NX4 MULT_OUT[3] NX154 NX233 MUX21_NI
        X_IX53 M_OUT_0 ADD_SIG MULT_OUT[4] NX52 MUX21_NI
        X_IX224 NX24 MULT_OUT[4] NX144 NX223 MUX21_NI
        X_IX214 NX24 MULT_OUT[5] NX134 NX213 MUX21_NI
*
.end
