* Component: /home/max/301/ECSE301_lab3/TopModel_S/TopModel  Viewpoint: ami05a
.OPTION VOLTAGE_LOOP_SEVERITY = WARNING
.INCLUDE /home/max/301/ECSE301_lab3/TopModel_S/TopModel/ami05a/TopModel_ami05a.spi
.INCLUDE /mgc/adk3_1/technology/ic/models/VDD_5.mod
.INCLUDE /mgc/adk3_1/technology/ic/models/ami05.mod
.PROBE TRAN V(DONE)
.PROBE TRAN V(MULT_OUT[0]) V(MULT_OUT[1]) V(MULT_OUT[2]) V(MULT_OUT[3])
+ V(MULT_OUT[4]) V(MULT_OUT[5]) V(MULT_OUT[6]) V(MULT_OUT[7])

VFORCE__Q_IN_2 Q_IN[2] GND dc 5

VFORCE__Q_IN_2_1_0 Q_IN[0] GND dc 0
VFORCE__Q_IN_2_1_1 Q_IN[1] GND dc
+ 0
VFORCE__Q_IN_2_1_2 Q_IN[3] GND dc 0

VFORCE__M_IN_0_0 M_IN[0] GND dc 5
VFORCE__M_IN_0_1 M_IN[1] GND dc 5

VFORCE__M_IN_2_0 M_IN[2] GND dc 0
VFORCE__M_IN_2_1 M_IN[3] GND dc 0

Vclock_0 CLOCK GND pattern 5 0 0 1n 1n 10n 0101 R
Vclock_1 CLOCK GND pattern 5 0
+ 0 1n 1n 10n 0101 R

VFORCE__START_0 START GND pattern 5 0 0 1n 1n 10n 1100
VFORCE__START_1 START GND
+ pattern 5 0 0 1n 1n 10n 1100




.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

.TEMP 27 

.TRAN  0 3000N 0 
